PLL4X_inst : PLL4X PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		c1	 => c1_sig,
		e0	 => e0_sig
	);
